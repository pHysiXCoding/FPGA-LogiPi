`timescale 1ns / 1ps

module main(
	iCLK_50,
			
	LED,
	PB,
	SW

   );
	input iCLK_50;

	input [1:0] LED;
	input [1:0] PB;
	input [1:0] SW;

	
	
	

endmodule
